module register_file (
    input clk,
    input rst,
    input write_enable,
    input  [4:0] rs1,
    input  [4:0] rs2, // add missing comma
    input  [4:0] rd1,
    input  [31:0] data_in,
    output [31:0] data1_out,
    output [31:0] data2_out
);

reg  [31:0] register [31:0];
integer i; // declare loop variable

// Register write part
always @(posedge clk) begin
    if (!rst) begin
        for (i  = 0; i < 32; i = i+1) begin
            register[i] <= 32'd0;
        end
    end else begin
        if (write_enable && (rd1 != 5'b0)) begin
            register[rd1] <= data_in;
        end
    end
end

assign data1_out = register[rs1];
assign data2_out = register[rs2]; 
endmodule